/*     Tambasis Georgios, aem 1797
	Axelos Christos, aem 1814
----------------------------------------
			
/*
  -to arxiko module
		-cpu-			
	-control_unit  + data_path-	 
 ------------ LIBRARY -----------
*/
`include "constants.h"

module CPU (clock, reset);
	input clock, reset;
	dataPath_controlUnit dataPath_controlUnit_0();
endmodule

	

	